library verilog;
use verilog.vl_types.all;
entity env_pkg is
end env_pkg;
