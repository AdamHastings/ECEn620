library verilog;
use verilog.vl_types.all;
entity my_package is
end my_package;
