library verilog;
use verilog.vl_types.all;
entity CovPort_pkg is
end CovPort_pkg;
