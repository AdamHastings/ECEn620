library verilog;
use verilog.vl_types.all;
entity transaction_pkg is
end transaction_pkg;
