library verilog;
use verilog.vl_types.all;
entity Driver_pkg is
end Driver_pkg;
