library verilog;
use verilog.vl_types.all;
entity Transaction_pkg is
end Transaction_pkg;
