library verilog;
use verilog.vl_types.all;
entity golden_module is
end golden_module;
