interface risc_spm_iface (input bit clk);

endinterface