library verilog;
use verilog.vl_types.all;
entity opcodes_include_v_unit is
end opcodes_include_v_unit;
