library verilog;
use verilog.vl_types.all;
entity ahb_if is
    port(
        clk             : in     vl_logic
    );
end ahb_if;
