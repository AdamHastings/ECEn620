library verilog;
use verilog.vl_types.all;
entity sram_if is
    port(
        clk             : in     vl_logic
    );
end sram_if;
