library verilog;
use verilog.vl_types.all;
entity arb_if is
    port(
        clk             : in     vl_logic
    );
end arb_if;
