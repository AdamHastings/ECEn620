library verilog;
use verilog.vl_types.all;
entity my_mem_if is
    port(
        clk             : in     vl_logic
    );
end my_mem_if;
