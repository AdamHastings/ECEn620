library verilog;
use verilog.vl_types.all;
entity Agent_pkg is
end Agent_pkg;
