library verilog;
use verilog.vl_types.all;
entity test is
    port(
        reset           : out    vl_logic
    );
end test;
