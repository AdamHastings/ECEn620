library verilog;
use verilog.vl_types.all;
entity Generator_pkg is
end Generator_pkg;
