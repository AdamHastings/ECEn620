library verilog;
use verilog.vl_types.all;
entity risc_spm_iface is
    port(
        clk             : in     vl_logic
    );
end risc_spm_iface;
